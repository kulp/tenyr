store[32'h00000000 + BASE] = 32'h41002004;
store[32'h00000001 + BASE] = 32'h42002005;
store[32'h00000002 + BASE] = 32'h03122006;
store[32'h00000003 + BASE] = 32'h00000000;
store[32'h00000004 + BASE] = 32'h73002123;
store[32'h00000005 + BASE] = 32'hffffffff;

`include "common.vh"
`timescale 1ms/10us

module lookup7(char, out);
    input[7:0] char;
    output reg[7:0] out = 0;

    always @(char) begin
        case (char)
           8'd032 /* ' ' */: out = 8'b11111111;
           8'd045 /* '-' */: out = 8'b10111111;

           8'd048 /* '0' */: out = 8'b11000000;
           8'd049 /* '1' */: out = 8'b11111001;
           8'd050 /* '2' */: out = 8'b10100100;
           8'd051 /* '3' */: out = 8'b10110000;
           8'd052 /* '4' */: out = 8'b10011001;
           8'd053 /* '5' */: out = 8'b10010010;
           8'd054 /* '6' */: out = 8'b10000010;
           8'd055 /* '7' */: out = 8'b11111000;
           8'd056 /* '8' */: out = 8'b10000000;
           8'd057 /* '9' */: out = 8'b10010000;

           8'd065 /* 'A' */: out = 8'b10001000;
           8'd067 /* 'C' */: out = 8'b11000110;
           8'd069 /* 'E' */: out = 8'b10000110;
           8'd070 /* 'F' */: out = 8'b10001110;
           8'd071 /* 'G' */: out = 8'b10000010;
           8'd072 /* 'H' */: out = 8'b10001001;
           8'd073 /* 'I' */: out = 8'b11111001;
           8'd074 /* 'J' */: out = 8'b11110001;
           8'd076 /* 'L' */: out = 8'b11000111;
           8'd079 /* 'O' */: out = 8'b11000000;
           8'd080 /* 'P' */: out = 8'b10001100;
           8'd083 /* 'S' */: out = 8'b10010010;
           8'd085 /* 'U' */: out = 8'b11000001;
           8'd089 /* 'Y' */: out = 8'b10010001;
           8'd090 /* 'Z' */: out = 8'b10100100;

           8'd098 /* 'b' */: out = 8'b10000011;
           8'd099 /* 'c' */: out = 8'b10100111;
           8'd100 /* 'd' */: out = 8'b10100001;
           8'd102 /* 'f' */: out = 8'b10001110;
           8'd103 /* 'g' */: out = 8'b10010000;
           8'd104 /* 'h' */: out = 8'b10001011;
           8'd105 /* 'i' */: out = 8'b11111001;
           8'd106 /* 'j' */: out = 8'b11110001;
           8'd111 /* 'o' */: out = 8'b10100011;
           8'd114 /* 'r' */: out = 8'b11100111;
           8'd117 /* 'u' */: out = 8'b11100011;
           8'd121 /* 'y' */: out = 8'b10010001;
           8'd122 /* 'z' */: out = 8'b10100100;

           default         : out = 8'b0xxxxxxx; // indicate bad digit with decimal point
        endcase
    end

endmodule


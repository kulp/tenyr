`include "common.vh"
`timescale 1ns/10ps

// External Interrupt Block
// contains its own RAMs and presents a simple interrupt handler interface
// to the tenyr Core
module Eib(input clk, reset_n, strobe, rw,
           input[IRQ_COUNT-1:0] irq, output reg trap,
           input[31:0] i_addr, output [31:0] i_data,
           input[31:0] d_addr, inout  [31:0] d_data);

    localparam IRQ_COUNT    = 32;               // total count of interrupts
    localparam DEPTH_BITS   = 2;                // maximum depth of stacks
    localparam MAX_DEPTH    = 1 << DEPTH_BITS;  // depth of stacks in words

    parameter  VEC_BOTTOM   = `VECTOR_ADDR;
    localparam VEC_BITS     = 5;                // vector table size in bits
    localparam VEC_SIZE     = 1 << VEC_BITS;    // vector table size in words
    parameter  VECTORFILE   = "vectors.memh";

    parameter  STACK_TOP    = `ISTACK_TOP;
    parameter  STACK_BITS   = 5;                // interrupt stack size in bits
    localparam STACK_SIZE   = 1 << STACK_BITS;  // interrupt stack size in words
    localparam STACK_WORDS  = (MAX_DEPTH << STACK_BITS) - 1;

    parameter  TRAMP_BOTTOM = `TRAMP_BOTTOM;
    parameter  TRAMP_BITS   = 6;                // trampoline size in bits
    localparam TRAMP_SIZE   = 1 << TRAMP_BITS;  // trampoline size in words

    // TODO use multidimensional array when tools support them
    //reg [31:0] stacks[STACK_WORDS:0];           // HW stack of interrupt stacks
    //reg [31:0] tramp[TRAMP_SIZE-1:0];           // single interrupt trampoline
    //reg [31:0] vecs[VEC_SIZE-1:0];              // interrupt vector table
    reg [31:0] rdata, i_rdata;                  // output on bus data lines
    //reg [31:0] stack_rdata, tramp_rdata, vecs_rdata;
    reg [31:0] stack_i_rdata, tramp_i_rdata, vecs_i_rdata;
    reg [31:0] stack_d_rdata, tramp_d_rdata, vecs_d_rdata;
    reg [31:0] stack_d_addr, tramp_d_addr, vecs_d_addr;
    reg [31:0] stack_i_addr, tramp_i_addr, vecs_i_addr;

    reg [DEPTH_BITS-1:0] depth = 0;             // stack pointer
    reg [ IRQ_COUNT-1:0] isr = 0;               // Interrupt Status Register
    reg [ IRQ_COUNT-1:0] imrs[MAX_DEPTH-1:0];   // Interrupt Mask Register stack
    reg [ IRQ_COUNT-1:0] rets[MAX_DEPTH-1:0];   // Return Address stack

    wire d_inrange = d_addr[31:12] == 20'hfffff;
    wire i_inrange = i_addr[31:12] == 20'hfffff;
    wire d_active  = d_inrange && strobe;
    assign d_data  = (d_active & ~rw) ? rdata : 32'bz;
    assign i_data  = i_inrange ? i_rdata : 32'bz;

    initial begin
        imrs[0] = 0;
        //$readmemh("../verilog/trampoline.memh", tramp.wrapped.store);
        //$readmemh(VECTORFILE, vecs.wrapped.store);
    end

`define IS_STACK(X)     ((STACK_TOP - STACK_SIZE) < (X) && (X) <= STACK_TOP)
`define IS_TRAMP(X)     (TRAMP_BOTTOM <= (X) && (X) < TRAMP_BOTTOM + TRAMP_SIZE)
`define IS_VEC(X)       (  VEC_BOTTOM <= (X) && (X) <   VEC_BOTTOM +   VEC_SIZE)
`define STACK_ADDR(X)   ((depth << STACK_BITS) | X[(STACK_BITS - 1):0])
`define TRAMP_ADDR(X)   (X[(TRAMP_BITS - 1):0])
`define VEC_ADDR(X)     (X[(VEC_BITS - 1):0])

    wire [31:0] vec_dout_d, vec_dout_i;
    wire [31:0] stack_dout_d, stack_dout_i;
    wire [31:0] tramp_dout_d, tramp_dout_i;

    wire [31:0]   vec_ad =   `VEC_ADDR(d_addr),   vec_ai =   `VEC_ADDR(i_addr);
    wire [31:0] stack_ad = `STACK_ADDR(d_addr), stack_ai = `STACK_ADDR(i_addr);
    wire [31:0] tramp_ad = `TRAMP_ADDR(d_addr), tramp_ai = `TRAMP_ADDR(i_addr);

    wire d_is_vec   = d_active && `IS_VEC  (d_addr), i_is_vec   = i_inrange && `IS_VEC  (i_addr);
    wire d_is_tramp = d_active && `IS_TRAMP(d_addr), i_is_tramp = i_inrange && `IS_TRAMP(i_addr);
    wire d_is_stack = d_active && `IS_STACK(d_addr), i_is_stack = i_inrange && `IS_STACK(i_addr);

    ramwrap #( // TODO vecs doesn't need to be accessible to instruction port
        .LOAD(1), .LOADFILE(VECTORFILE), .ABITS(VEC_BITS), .SIZE(VEC_SIZE)
    ) vecs(
        .clka  ( clk            ), .clkb  ( clk        ),
        .ena   ( d_is_vec       ), .enb   ( i_is_vec   ),
        .wea   ( d_active && rw ), .web   ( 1'b0       ),
        .addra ( vec_ad         ), .addrb ( vec_ai     ),
        .dina  ( d_data         ), .dinb  ( 32'bx      ),
        .douta ( vec_dout_d     ), .doutb ( vec_dout_i )
    );

    ramwrap #(.ABITS(STACK_BITS), .SIZE(STACK_SIZE)) stack(
        .clka  ( clk            ), .clkb  ( clk          ),
        .ena   ( d_is_stack     ), .enb   ( i_is_stack   ),
        .wea   ( d_active && rw ), .web   ( 1'b0         ),
        .addra ( stack_ad       ), .addrb ( stack_ai     ),
        .dina  ( d_data         ), .dinb  ( 32'bx        ),
        .douta ( stack_dout_d   ), .doutb ( stack_dout_i )
    );

    ramwrap #(.ABITS(TRAMP_BITS), .SIZE(TRAMP_SIZE)) tramp(
        .clka  ( clk            ), .clkb  ( clk          ),
        .ena   ( d_is_tramp     ), .enb   ( i_is_tramp   ),
        .wea   ( d_active && rw ), .web   ( 1'b0         ),
        .addra ( tramp_ad       ), .addrb ( tramp_ai     ),
        .dina  ( d_data         ), .dinb  ( 32'bx        ),
        .douta ( tramp_dout_d   ), .doutb ( tramp_dout_i )
    );

    always @(posedge clk) begin
        if (!reset_n) begin
            isr     <= 0;
            depth   <= 0;
            imrs[0] <= 0;
        end else begin
            isr  <= isr | irq;  // accumulate until cleared
            // For now, trap follows irq by one cycle
            trap <= |(imrs[depth] & isr);

            if (d_active && rw) begin // writing
                if (!(d_is_vec | d_is_tramp | d_is_stack)) case (d_addr[11:0])
                    12'hfff: begin
                        if (depth == MAX_DEPTH - 1) begin
                            $display("Tried to push too many interrupt frames");
                            $stop;
                        end else
                            depth <= depth + 1;

                        rets[depth + 1] <= d_data;
                        imrs[depth + 1] <= 'b0;     // disable interrupts
                    end
                    12'hffe: isr <= isr & ~d_data;    // ISR clear bits
                    12'hffd: imrs[depth] <= d_data;   // IMR write
                    default: $display("Unhandled write of %x @ %x", d_data, d_addr);
                endcase
            end else if (d_inrange) begin   // reading
                     if (d_is_stack) rdata <= stack_dout_d;
                else if (d_is_tramp) rdata <= tramp_dout_d;
                else if (d_is_vec  ) rdata <= vec_dout_d;
                else case (d_addr[11:0])
                    12'hfff: begin
                        if (d_active) begin
                            if (depth == 0) begin
                                $display("Tried to pop too many interrupt frames");
                                $stop;
                            end else
                                depth <= depth - 1;
                        end

                        rdata <= rets[depth];       // RA  read
                    end
                    12'hffe: rdata <= isr;          // ISR read
                    12'hffd: rdata <= imrs[depth];  // IMR read
                    default: if (d_active) $display("Unhandled read @ %x", d_addr);
                endcase
            end
        end
    end

endmodule


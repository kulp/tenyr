`include "common.vh"
`timescale 1ms/10us

module lookup7(input[7:0] char, output[6:0] lines);
    reg[6:0] out = 7'b0;
    assign lines = out;

    case (char)
       8'd045 /* '-' */: out = 7'b0000001;

       8'd065 /* 'A' */: out = 7'b1110111;
       8'd067 /* 'C' */: out = 7'b1001110;
       8'd069 /* 'E' */: out = 7'b1001111;
       8'd070 /* 'F' */: out = 7'b1000111;
       8'd071 /* 'G' */: out = 7'b1011111;
       8'd072 /* 'H' */: out = 7'b0110111;
       8'd073 /* 'I' */: out = 7'b0110000;
       8'd074 /* 'J' */: out = 7'b0111000;
       8'd076 /* 'L' */: out = 7'b0001110;
       8'd079 /* 'O' */: out = 7'b1111110;
       8'd080 /* 'P' */: out = 7'b1100111;
       8'd083 /* 'S' */: out = 7'b1011011;
       8'd085 /* 'U' */: out = 7'b0111110;
       8'd089 /* 'Y' */: out = 7'b0111011;
       8'd090 /* 'Z' */: out = 7'b1101101;

       8'd098 /* 'b' */: out = 7'b0011111;
       8'd099 /* 'c' */: out = 7'b0001101;
       8'd100 /* 'd' */: out = 7'b0111101;
       8'd102 /* 'f' */: out = 7'b1000111;
       8'd103 /* 'g' */: out = 7'b1111011;
       8'd104 /* 'h' */: out = 7'b0010111;
       8'd105 /* 'i' */: out = 7'b0110000;
       8'd106 /* 'j' */: out = 7'b0111000;
       8'd111 /* 'o' */: out = 7'b0011101;
       8'd117 /* 'u' */: out = 7'b0011100;
       8'd121 /* 'y' */: out = 7'b0111011;
       8'd122 /* 'z' */: out = 7'b1101101;

       8'd048 /* '0' */: out = 7'b1111110;
       8'd049 /* '1' */: out = 7'b0110000;
       8'd050 /* '2' */: out = 7'b1101101;
       8'd051 /* '3' */: out = 7'b1111001;
       8'd052 /* '4' */: out = 7'b0110011;
       8'd053 /* '5' */: out = 7'b1011011;
       8'd054 /* '6' */: out = 7'b1011111;
       8'd055 /* '7' */: out = 7'b1110000;
       8'd056 /* '8' */: out = 7'b1111111;
       8'd057 /* '9' */: out = 7'b1111011;
    endcase

endmodule

